// 라운드 끝나고 matchresult랑 클럭 입력되면
// round counter, win counter, lose counter 업데이트

// Lab6에 counter 모듈 쓰기

// round는 라운드 끝날때마다 1 추가
// p1 승이면 win counter 1 추가
// p2 승이면 lose counter 1 추가

module counter(
    

);

endmodule